module breath_led(
    input          sys_clk        , //??????
    input          sys_rst_n      , //??????
    input          sw_ctrl        , //??????????????? 1???? 0:??
    input          set_en         , //??????????????????????
    input   [9:0]  set_freq_step  , //????????????c????
    
    output         led              //LED
);

//*****************************************************
//**                  main code
//*****************************************************

//parameter define
parameter  START_FREQ_STEP = 10'd100; //??????????????

//reg define
reg  [15:0]  period_cnt  ;      //?????????
reg  [9:0]   freq_step   ;      //???????????????
reg  [15:0]  duty_cycle  ;      //?????????????????
reg          inc_dec_flag;      //???????????????????,???????????
                                //?1??????????,?0???????????
//wire define
wire         led_t       ;


assign led_t = ( period_cnt <= duty_cycle ) ? 1'b1 : 1'b0 ;
assign led = led_t & sw_ctrl;

//??????????????0-50_000??????
always @ (posedge sys_clk) begin
    if (!sys_rst_n)
        period_cnt <= 16'd0;
    else if(!sw_ctrl)
        period_cnt <= 16'd0;
    else if( period_cnt == 16'd50_000 )
        period_cnt <= 16'd0;
    else
        period_cnt <= period_cnt + 16'd1;
end

//?????????
always @(posedge sys_clk) begin
    if(!sys_rst_n)
        freq_step <= START_FREQ_STEP;
    else if(set_en) begin
        if(set_freq_step == 0)
            freq_step <= 10'd1;
        else if(set_freq_step >= 10'd1_000)
            freq_step <= 10'd1_000;
        else    
            freq_step <= set_freq_step;
    end        
end

//???????????????
always @(posedge sys_clk) begin
    if (sys_rst_n == 1'b0) begin
        duty_cycle <= 16'd0;
        inc_dec_flag <= 1'b0;
    end     
    else if(!sw_ctrl) begin          //?????????????????????
        duty_cycle <= 16'd0;
        inc_dec_flag <= 1'b0;
    end    
    //???????????????????????????????
    else if( period_cnt == 16'd50_000 ) begin
        if( inc_dec_flag ) begin  //??????
            if( duty_cycle == 16'd0 )     
                inc_dec_flag <= 1'b0;
            else if(duty_cycle < freq_step)
                duty_cycle <= 16'd0;
            else    
                duty_cycle <= duty_cycle - freq_step;
        end
        else begin  //???????
            if( duty_cycle >= 16'd50_000 )  
                inc_dec_flag <= 1'b1;
            else
                duty_cycle <= duty_cycle + freq_step;
        end 
    end 
    else  //???????????????????????????
        duty_cycle <= duty_cycle ;
end
  
endmodule